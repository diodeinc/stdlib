V1 VCC GND SIN(0 5V 1kHz)

.control
  tran 0.01m 5m
  plot v(VCC) v(PROBE)
.endc
