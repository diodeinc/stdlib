V1 VCC GND SIN(0 5V 1kHz)

.control
  tran 0.001m 5m
  plot v(VCC) v(PROBE)
  
  * Save the output to 
  set hcopydevtype = svg
  hardcopy build/sim.svg v(VCC) v(PROBE)
  quit
.endc
